`define CODE 12'h000
`define DATA 12'h001
`define VGA  12'h002
`define KBD  12'h003
`define LED  12'h004
`define HEX  12'h005
`define CLK  12'h006
`define SW   12'h007